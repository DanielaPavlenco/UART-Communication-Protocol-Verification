  // Add necessary interface signals and methods
  // Example: tx, rx, baud_rate, etc.

  // Add your interface logic here

endinterface : UART_Interface
